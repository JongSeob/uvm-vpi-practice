// Code your testbench here
// or browse Examples
module tb;
  
  initial begin
    $display("Hello Questa!\n");
    $hello();
  end
  
endmodule